--Steven Miller
--11710
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use ieee.NUMERIC_STD.UNSIGNED;

entity rom_tb is
end rom_tb;

architecture TB of rom_tb is
component ROM is
PORT
(
	address		: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
	clock		: IN STD_LOGIC  := '1';
	rden		: IN STD_LOGIC  := '1';
	q		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
);
end component;

signal address : std_logic_vector(9 downto 0);
signal clock : std_logic;
signal rden : std_logic;
signal q : std_logic_vector(31 downto 0);
begin  -- TB

  UUT : ROM
    port map 
(
      --inputs => inputs,
      clock    => clock,
      q => q,
      address => address,
      rden=>rden
      
);

clock <= not(clock) after 10 ns;

process

--wait for 10ns
--check output

begin
--wait for filter to start up
--resetn<='1';
rden <= '1';
for i in 0 to 1023 loop
	address <= STD_LOGIC_VECTOR(to_unsigned(i,address'length));
	wait until rising_edge(clock);
	end loop;

end process;
end TB;